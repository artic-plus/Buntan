module inv_test(A,Y);
    input A;
    output Y;
    assign Y = !A;
endmodule